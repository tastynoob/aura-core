`include "backend_define.svh"






module dcache #(
    parameter int BANKS = 4,
    parameter int SETS = 4,
    parameter int WAYS = 4,
    parameter int ADDRWIDTH = `PALEN,
    parameter int CACHELINSIZE = `CACHELINE_SIZE
) (

);






endmodule


