
module tb (
    input clk,
    input rst
);

`ifdef DEBUG
// refcount u_refcount(
//     .clk                  (clk                  ),
//     .rst                  (rst                  ),
//     .i_alloc_ismv         (         ),
//     .i_alloc_req          (          ),
//     .i_alloc_prIdx        (        ),
//     .i_dealloc_req        (        ),
//     .i_dealloc_prIdx      (      ),
//     .o_real_dealloc_req   (   ),
//     .o_real_dealloc_prIdx ( )
// );

`endif

endmodule


