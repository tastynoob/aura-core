
`include "core_define.svh"

module tb (
    input clk,
    input rst
);

`ifdef DEBUG




`endif

endmodule




