`ifndef __CORE_SPEC_SVH__
`define __CORE_SPEC_SVH__


`define SV39_SUPPORT 1

`define PALEN 36

`define VADDR(x) ``x``[39-1:0]











`endif
