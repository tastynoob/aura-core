



interface issueport_if;




endinterface
