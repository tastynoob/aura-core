


module rob();

endmodule
