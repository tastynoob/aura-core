


module ROB();

endmodule
