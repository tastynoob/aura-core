
`include "core_define.svh"
`include "frontend_define.svh"

module tb (
    input wire clk,
    input wire rst
);





endmodule



