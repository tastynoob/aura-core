




// cpu frontend
// storage <-tilelink-> frontend <--> backend




module aura_frontend (
    input wire clk,
    input wire rst,


    // to next level storage
    tilelink_if.m if_fetch_bus
);









endmodule



