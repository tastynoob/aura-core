`ifndef __DISPATCH_DEFINE_SVH__
`define __DISPATCH_DEFINE_SVH__

`include "core_define.svh"


// TODO: we may need to implement pcbuffer and immbuffer

//dispatch queue type
`define DQ_INT 0
`define DQ_MEM 1






`endif
