`include "dispatch_define.svh"




module dispQue #(
    parameter int DEPTH = 4,
    parameter int INPORT_NUM  = `RENAME_WIDTH,
    parameter int OUTPORT_NUM = 4,
    parameter int DQTYPE = 0
) (
    input wire clk,
    input wire rst
);










endmodule








